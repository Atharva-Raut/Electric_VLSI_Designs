*** SPICE deck for cell Two_Stage_OTA{lay} from library Amplifiers
*** Created on Sat Jul 17, 2021 00:44:12
*** Last revised on Sun Jul 18, 2021 00:56:17
*** Written on Sun Jul 18, 2021 00:56:24 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: Two_Stage_OTA{lay}
Mnmos@0 net@1 V_out net@0 gnd nMOS L=0.6U W=3.6U AS=7.02P AD=5.783P PS=11.1U PD=7.2U
Mnmos@1 net@3 V+ net@1 gnd nMOS L=0.6U W=3.6U AS=5.783P AD=7.02P PS=7.2U PD=11.1U
Mnmos@2 net@1 V_b gnd gnd nMOS L=0.6U W=3.6U AS=14.22P AD=5.783P PS=21.7U PD=7.2U
Mnmos@3 gnd V_b net@1 gnd nMOS L=0.6U W=3.6U AS=5.783P AD=14.22P PS=7.2U PD=21.7U
Mnmos@4 V_out V_b gnd gnd nMOS L=0.6U W=3.6U AS=14.22P AD=7.02P PS=21.7U PD=11.1U
Mpmos@0 vdd net@0 net@0 vdd pMOS L=0.6U W=3.6U AS=7.02P AD=12.42P PS=11.1U PD=18.3U
Mpmos@1 net@3 net@0 vdd vdd pMOS L=0.6U W=3.6U AS=12.42P AD=7.02P PS=18.3U PD=11.1U
Mpmos@2 V_out net@3 vdd vdd pMOS L=0.6U W=3.6U AS=12.42P AD=7.02P PS=18.3U PD=11.1U

* Spice Code nodes in cell cell 'Two_Stage_OTA{lay}'
vdd VDD 0 DC 5
vin V+ 0 pulse(0 5 0 1us 0)
vin2 V_b 0 DC 1.0
.tran 1us
.include C:\Users\athar\Documents\Electric VLSI\C5_models.txt
.END
